# ====================================================================
#
#      flash_intel_28fxxx.cdl
#
#      FLASH memory - Hardware support for Intel flash parts
#
# ====================================================================
### ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2009 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Contributors:   jskov, gthomas
# Date:           2001-03-21
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_INTEL_28FXXX {
    display       "Intel FlashFile FLASH memory support"
    description   "FLASH memory device support for Intel FlashFile"
    parent        CYGPKG_IO_FLASH
    active_if	  CYGPKG_IO_FLASH

    active_if     CYGINT_DEVS_FLASH_INTEL_28FXXX_REQUIRED

    implements    CYGHWR_IO_FLASH_DEVICE
    implements    CYGHWR_IO_FLASH_DEVICE_LEGACY

    include_dir   cyg/io

    requires      { CYGINT_DEVS_FLASH_INTEL_VARIANTS != 0 }

    cdl_option CYGNUM_DEVS_FLASH_INTEL_28FXXX_TIMEOUT {
        display       "Timeout for flash operations (simple counter based)"
        flavor        data
        legal_values  1000000 to 1000000000
        default_value 50000000
        description   " 
            Timeout for flash operations. This is just a simple
            counter. It depends on the speed of the flash, the processor, etc.
            It has to be adjusted for each hardware configuration. "
    }


    cdl_interface CYGINT_DEVS_FLASH_INTEL_VARIANTS {
        display   "Number of included variants"
    }

    cdl_interface CYGHWR_DEVS_FLASH_INTEL_BUFFERED_WRITES {
        flavor    booldata
        display   "Must support buffered writes"
    }

    cdl_option CYGHWR_DEVS_FLASH_INTEL_28F160S5 {
        display       "Intel 28F160S5 flash memory support"
        default_value 0
        implements    CYGINT_DEVS_FLASH_INTEL_VARIANTS
        implements    CYGHWR_DEVS_FLASH_INTEL_BUFFERED_WRITES
        description   "
            When this option is enabled, the Intel flash driver will be
            able to recognize and handle the 28F160S5
            part in the family."
    }

    cdl_option CYGHWR_DEVS_FLASH_INTEL_28F160B3T {
        display       "Intel 28F160B3T flash memory support"
        default_value 0
        implements    CYGHWR_IO_FLASH_BLOCK_LOCKING
        implements    CYGINT_DEVS_FLASH_INTEL_VARIANTS
        description   "
            When this option is enabled, the Intel flash driver will be
            able to recognize and handle the 28F160B3T
            part in the family."
    }

    cdl_option CYGHWR_DEVS_FLASH_INTEL_28F160C3B {
        display       "Intel 28F160C3B flash memory support"
        default_value 0
        implements    CYGHWR_IO_FLASH_BLOCK_LOCKING
        implements    CYGINT_DEVS_FLASH_INTEL_VARIANTS
        description   "
            When this option is enabled, the Intel flash driver will be
            able to recognize and handle the 28F160C3B
            part in the family."
    }

    cdl_option CYGHWR_DEVS_FLASH_INTEL_28F320B3 {
        display       "Intel 28F320B3 flash memory support"
        default_value 0
        implements    CYGINT_DEVS_FLASH_INTEL_VARIANTS
        description   "
            When this option is enabled, the Intel flash driver will be
            able to recognize and handle the 28F320B3
            part in the family."
    }


    cdl_option CYGHWR_DEVS_FLASH_INTEL_28F320C3 {
        display       "Intel 28F320C3 flash memory support"
        default_value 0
        implements    CYGHWR_IO_FLASH_BLOCK_LOCKING
        implements    CYGINT_DEVS_FLASH_INTEL_VARIANTS
        description   "
            When this option is enabled, the Intel flash driver will be
            able to recognize and handle the 28F320C3
            part in the family."
    }

    cdl_option CYGHWR_DEVS_FLASH_INTEL_28F320S3 {
        display       "Intel 28F320S3 flash memory support"
        default_value 0
        implements    CYGHWR_IO_FLASH_BLOCK_LOCKING
        implements    CYGINT_DEVS_FLASH_INTEL_VARIANTS
        description   "
            When this option is enabled, the Intel flash driver will be
            able to recognize and handle the 28F320S3
            part in the family."
    }

    cdl_option CYGHWR_DEVS_FLASH_INTEL_28F128K3 {
        display       "Intel 28F128K3 flash memory support"
        default_value 0
        implements    CYGHWR_IO_FLASH_BLOCK_LOCKING
        implements    CYGINT_DEVS_FLASH_INTEL_VARIANTS
        description   "
            When this option is enabled, the Intel flash driver will be
            able to recognize and handle the 28F128K3
            part in the family."
    }

   cdl_option CYGHWR_DEVS_FLASH_INTEL_28F128P30 {
        display       "Intel 28F128P30 flash memory support"
        default_value 0
        implements    CYGHWR_IO_FLASH_BLOCK_LOCKING
        implements    CYGINT_DEVS_FLASH_INTEL_VARIANTS
        implements    CYGHWR_DEVS_FLASH_INTEL_BUFFERED_WRITES
        description   "
            When this option is enabled, the Intel flash driver will be
            able to recognize and handle the 28F128P30
            part in the family."
    }

    cdl_option CYGHWR_DEVS_FLASH_INTEL_28F128J3 {
        display       "Intel 28F128J3 flash memory support"
        default_value 0
        implements    CYGHWR_IO_FLASH_BLOCK_LOCKING
        implements    CYGINT_DEVS_FLASH_INTEL_VARIANTS
        description   "
            When this option is enabled, the Intel flash driver will be
            able to recognize and handle the 28F128J3
            part in the family."
    }

    cdl_option CYGHWR_DEVS_FLASH_INTEL_28F320J3 {
        display       "Intel 28F320J3 flash memory support"
        default_value 0
        implements    CYGHWR_IO_FLASH_BLOCK_LOCKING
        implements    CYGINT_DEVS_FLASH_INTEL_VARIANTS
        description   "
            When this option is enabled, the Intel flash driver will be
            able to recognize and handle the 28F320J3
            part in the family."
    }

    cdl_option CYGHWR_DEVS_FLASH_INTEL_28F800B5 {
        display       "Intel 28F800B5 flash memory support"
        default_value 0
        implements    CYGINT_DEVS_FLASH_INTEL_VARIANTS
        description   "
            When this option is enabled, the Intel flash driver will be
            able to recognize and handle the 28F800B5
            part in the family."
    }

    cdl_option CYGHWR_DEVS_FLASH_SHARP_LH28F016SCT_Z4 {
        display       "Sharp LH28F016SCT-Z4 flash memory support"
        default_value 0
        implements    CYGHWR_IO_FLASH_BLOCK_LOCKING
        implements    CYGINT_DEVS_FLASH_INTEL_VARIANTS
        description   "
            When this option is enabled, the Intel flash driver will be
            able to recognize and handle the Sharp LH28F016SCT-Z4
            part.  Although this part is not an Intel part, the driver
            is implemented using the same command status definitions."

    }

    cdl_option CYGHWR_DEVS_FLASH_SHARP_LH28F016SCT_95 {
        display       "Sharp LH28F016SCT-95 flash memory support"
        default_value 0
        implements    CYGHWR_IO_FLASH_BLOCK_LOCKING
        implements    CYGINT_DEVS_FLASH_INTEL_VARIANTS
        description   "
            When this option is enabled, the Intel flash driver will be
            able to recognize and handle the Sharp LH28F016SCT-95
            part.  Although this part is not an Intel part, the driver
            is implemented using the same command status definitions."

    }
    cdl_option CYGHWR_DEVS_FLASH_INTEL_JS28F640P30B85 {
 		display       "Intel JS28F640P30B85 flash memory support"
        default_value 1
        implements    CYGHWR_IO_FLASH_BLOCK_LOCKING
        implements    CYGINT_DEVS_FLASH_INTEL_VARIANTS
        description   "
            When this option is enabled, the Intel flash driver will be
            able to recognize and handle the JS28F640P30B85
            part in the family."
    }
    
}
